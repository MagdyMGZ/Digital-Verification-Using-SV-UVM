package Wrapper_pack ;
	typedef enum bit[2:0] {IDLE,CHK_CMD,WRITE,READ_ADD,READ_DATA} state_e ;
endpackage 

